
module lab3_sys (
	clk_clk,
	i2c_scl_pad_io,
	i2c_sda_pad_io,
	pio_0_seg_export,
	pio_1_btn_export,
	reset_reset_n);	

	input		clk_clk;
	inout		i2c_scl_pad_io;
	inout		i2c_sda_pad_io;
	output	[23:0]	pio_0_seg_export;
	input		pio_1_btn_export;
	input		reset_reset_n;
endmodule
